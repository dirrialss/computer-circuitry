module ref_sum (Ain, Bin, Ci, Sout, Co);
  input [7:0] Ain, Bin;  // ????????? ??????????? ?? 8 ???
  input Ci;
  output [7:0] Sout;     // ????????? ??????????? ?? 8 ???
  output Co;
  reg [8:0] S;           // ????????? ??????????? ?? 9 ??? (8 ??? + ???????????)
  
  // ?????????? ???? ?? ????????????? ?????
  always @ (Ain or Bin or Ci)
    S = Ain + Bin + Ci;
    
  // ???????? ??????????: ??????? 8 ??? - ????, ??????? ??? - ???????????
  assign Sout = S[7:0];
  assign Co = S[8];
endmodule
