library verilog;
use verilog.vl_types.all;
entity multiplexer_8to1_tb is
end multiplexer_8to1_tb;
