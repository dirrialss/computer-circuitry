library verilog;
use verilog.vl_types.all;
entity comb2_Siukalo is
    port(
        x3              : in     vl_logic;
        x2              : in     vl_logic;
        x1              : in     vl_logic;
        f4              : out    vl_logic
    );
end comb2_Siukalo;
